`timescale 1ns/1ps
module tt_um_turbo_codec (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

    // Input/Output assignments
    wire data_in = ui_in[0];
    wire start = ui_in[1];
    wire encode_mode = ui_in[2];  // 1=encode, 0=decode
    wire reset = ~rst_n;
    
    // Output assignments
    assign uo_out[0] = encoded_out[0];
    assign uo_out[1] = encoded_out[1];
    assign uo_out[2] = encoded_out[2];
    assign uo_out[3] = decoded_out;
    assign uo_out[4] = output_valid;
    assign uo_out[7:5] = 3'b000;
    
    // Unused IOs
    assign uio_out = 8'b0;
    assign uio_oe = 8'b0;
    
    // Internal signals
    reg [2:0] encoded_out;
    reg decoded_out;
    reg output_valid;
    
    // Encoder signals
    wire [2:0] encoder_output;
    wire encoder_valid;
    
    // Decoder signals
    wire decoder_output;
    wire decoder_valid;
    
    // Select between encoder and decoder outputs
    always @(posedge clk) begin
        if (reset) begin
            encoded_out <= 3'b0;
            decoded_out <= 1'b0;
            output_valid <= 1'b0;
        end else begin
            if (encode_mode) begin
                encoded_out <= encoder_output;
                decoded_out <= 1'b0;
                output_valid <= encoder_valid;
            end else begin
                encoded_out <= 3'b0;
                decoded_out <= decoder_output;
                output_valid <= decoder_valid;
            end
        end
    end
    
    // Instantiate Turbo Encoder
    turbo_encoder encoder_inst (
        .clk(clk),
        .reset(reset),
        .data_in(data_in),
        .start(start & encode_mode),
        .encoded_out(encoder_output),
        .valid(encoder_valid)
    );
    
    // Instantiate Turbo Decoder
    turbo_decoder decoder_inst (
        .clk(clk),
        .reset(reset),
        .encoded_in({ui_in[5:3]}), // 3-bit encoded input
        .start(start & ~encode_mode),
        .decoded_out(decoder_output),
        .valid(decoder_valid)
    );

endmodule

// Turbo Encoder Module
module turbo_encoder (
    input wire clk,
    input wire reset,
    input wire data_in,
    input wire start,
    output reg [2:0] encoded_out,
    output reg valid
);

    // RSC (Recursive Systematic Convolutional) encoder parameters
    // Generator polynomials: G1 = 1+D+D^3, G2 = 1+D^2+D^3
    parameter G1 = 4'b1011; // 1+D+D^3
    parameter G2 = 4'b1101; // 1+D^2+D^3
    
    // State registers for two constituent encoders
    reg [2:0] state1, state2;
    reg [3:0] shift_reg1, shift_reg2;
    
    // Interleaver (simplified - fixed pattern for 8-bit block)
    reg [7:0] interleaver_pattern = 8'h45; // Simple pattern
    reg [2:0] bit_counter;
    reg [7:0] input_buffer;
    reg encoding_active;
    
    // Parity calculation functions
    function parity_calc;
        input [3:0] data;
        input [3:0] gen_poly;
        begin
            parity_calc = ^(data & gen_poly);
        end
    endfunction
    
    always @(posedge clk) begin
        if (reset) begin
            state1 <= 3'b0;
            state2 <= 3'b0;
            shift_reg1 <= 4'b0;
            shift_reg2 <= 4'b0;
            bit_counter <= 3'b0;
            input_buffer <= 8'b0;
            encoding_active <= 1'b0;
            encoded_out <= 3'b0;
            valid <= 1'b0;
        end else begin
            if (start && !encoding_active) begin
                encoding_active <= 1'b1;
                bit_counter <= 3'b0;
                input_buffer[bit_counter] <= data_in;
                valid <= 1'b0;
            end else if (encoding_active) begin
                if (bit_counter < 7) begin
                    bit_counter <= bit_counter + 1;
                    input_buffer[bit_counter + 1] <= data_in;
                end else begin
                    // Start encoding process
                    // Systematic bit
                    encoded_out[0] <= input_buffer[0];
                    
                    // First parity bit (encoder 1)
                    shift_reg1 <= {shift_reg1[2:0], input_buffer[0]};
                    encoded_out[1] <= parity_calc(shift_reg1, G1);
                    
                    // Second parity bit (encoder 2) - with interleaving
                    shift_reg2 <= {shift_reg2[2:0], input_buffer[interleaver_pattern[2:0]]};
                    encoded_out[2] <= parity_calc(shift_reg2, G2);
                    
                    valid <= 1'b1;
                    encoding_active <= 1'b0;
                end
            end else begin
                valid <= 1'b0;
            end
        end
    end

endmodule

// Turbo Decoder Module (Simplified BCJR Algorithm)
module turbo_decoder (
    input wire clk,
    input wire reset,
    input wire [2:0] encoded_in,
    input wire start,
    output reg decoded_out,
    output reg valid
);

    // Simplified decoder states
    reg [1:0] decoder_state;
    reg [3:0] iteration_count;
    reg decoding_active;
    
    // LLR (Log-Likelihood Ratio) storage (simplified)
    reg signed [7:0] llr_systematic;
    reg signed [7:0] llr_parity1;
    reg signed [7:0] llr_parity2;
    reg signed [7:0] extrinsic_info;
    
    // Decoder parameters
    parameter MAX_ITERATIONS = 4;
    parameter LLR_SCALE = 8; // Scaling factor for LLR values
    
    always @(posedge clk) begin
        if (reset) begin
            decoder_state <= 2'b00;
            iteration_count <= 4'b0;
            decoding_active <= 1'b0;
            decoded_out <= 1'b0;
            valid <= 1'b0;
            llr_systematic <= 8'b0;
            llr_parity1 <= 8'b0;
            llr_parity2 <= 8'b0;
            extrinsic_info <= 8'b0;
        end else begin
            case (decoder_state)
                2'b00: begin // Idle
                    if (start && !decoding_active) begin
                        decoding_active <= 1'b1;
                        decoder_state <= 2'b01;
                        iteration_count <= 4'b0;
                        
                        // Initialize LLRs based on received symbols
                        llr_systematic <= encoded_in[0] ? LLR_SCALE : -LLR_SCALE;
                        llr_parity1 <= encoded_in[1] ? LLR_SCALE : -LLR_SCALE;
                        llr_parity2 <= encoded_in[2] ? LLR_SCALE : -LLR_SCALE;
                        
                        valid <= 1'b0;
                    end
                end
                
                2'b01: begin // First decoder processing
                    // Simplified BCJR algorithm for first constituent decoder
                    extrinsic_info <= llr_systematic + llr_parity1;
                    decoder_state <= 2'b10;
                end
                
                2'b10: begin // Second decoder processing
                    // Simplified BCJR algorithm for second constituent decoder
                    extrinsic_info <= extrinsic_info + llr_parity2;
                    
                    if (iteration_count < MAX_ITERATIONS - 1) begin
                        iteration_count <= iteration_count + 1;
                        decoder_state <= 2'b01; // Go back for another iteration
                    end else begin
                        decoder_state <= 2'b11; // Final decision
                    end
                end
                
                2'b11: begin // Final decision and output
                    decoded_out <= (extrinsic_info > 0) ? 1'b1 : 1'b0;
                    valid <= 1'b1;
                    decoding_active <= 1'b0;
                    decoder_state <= 2'b00;
                end
                
                default: decoder_state <= 2'b00;
            endcase
        end
    end

endmodule

